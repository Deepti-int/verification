class a ;
  int data;
  but [7:0]addr;
endclass

