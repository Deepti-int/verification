class base;
  int data;
  bit[7:0]addr;
endclass

class child extends base;
endclass
